module divide_32(
	input [31:0] Ra, Rb,
	output [31:0] quotient, remainder
	);
	remainder = Ra%Rb;
	quoitent = (Ra-remainder)/Rb
	
endmodule