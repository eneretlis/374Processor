module c_flipflop(input D, C
						output Q);
	always @(posedge C)
	begin 
		Q <= D;
	end
endmodule
